-------------------------------------------------------------------------------
--   ____  ____ 
--  /   /\/   / 
-- /___/  \  /    Vendor: Xilinx 
-- \   \   \/     Version : 3.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard  
--  /   /         Filename : gtwizard_v2_5_gt_frame_check.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\ 
--
--
-- Module gtwizard_v2_5_GT_FRAME_CHECK
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard  
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;
use ieee.std_logic_textio.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

--***********************************Entity Declaration************************

entity gtwizard_v2_5_GT_FRAME_CHECK is
generic
(
    RX_DATA_WIDTH            : integer := 16;
    RXCTRL_WIDTH             : integer := 2;
    WORDS_IN_BRAM            : integer := 256;
    CHANBOND_SEQ_LEN         : integer := 1;
    COMMA_DOUBLE             : std_logic_vector(15 downto 0) := x"f628";
    START_OF_PACKET_CHAR     : std_logic_vector (15 downto 0)  := x"02bc"
);
port
(
    -- User Interface
    RX_DATA_IN               : in  std_logic_vector((RX_DATA_WIDTH-1) downto 0); 
    RXCTRL_IN                : in  std_logic_vector((RXCTRL_WIDTH-1) downto 0);

    RXENPCOMMADET_OUT        : out std_logic;
    RXENMCOMMADET_OUT        : out std_logic;
    RX_ENCHAN_SYNC_OUT       : out std_logic;
    RX_CHANBOND_SEQ_IN       : in  std_logic;

    -- Control Interface
    INC_IN                   : in  std_logic; 
    INC_OUT                  : out std_logic; 
    PATTERN_MATCHB_OUT       : out std_logic;
    RESET_ON_ERROR_IN        : in  std_logic;


    -- Error Monitoring
    ERROR_COUNT_OUT          : out std_logic_vector(7 downto 0);
    
    -- Track Data
    TRACK_DATA_OUT           : out std_logic;

    RX_SLIDE                  : out std_logic;
    -- System Interface
    USER_CLK                 : in std_logic;       
    SYSTEM_RESET             : in std_logic
  
);


end gtwizard_v2_5_GT_FRAME_CHECK;

architecture RTL of gtwizard_v2_5_GT_FRAME_CHECK is
    attribute DowngradeIPIdentifiedWarnings: string;
    attribute DowngradeIPIdentifiedWarnings of RTL : architecture is "yes";
--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

--***************************Internal Register Declarations********************
    signal  reset_on_error_in_r         :   std_logic;
    signal  reset_on_error_in_r2         :   std_logic;
    signal  system_reset_r              :   std_logic;
    signal  system_reset_r2              :   std_logic;
    attribute keep: string;
    attribute keep of system_reset_r    :   signal is "true";
    attribute keep of system_reset_r2    :   signal is "true";
    attribute ASYNC_REG                        : string;
     attribute ASYNC_REG of system_reset_r     : signal is "TRUE";
     attribute ASYNC_REG of system_reset_r2     : signal is "TRUE";

    signal  begin_r                     :   std_logic;
    signal  data_error_detected_r       :   std_logic;
    signal  error_count_r               :   unsigned(8 downto 0);
    signal  error_detected_r            :   std_logic;
    signal  read_counter_i              :   unsigned(9 downto 0);    
    signal  read_counter_conv           :   std_logic_vector(9 downto 0);    
    signal  rx_data_r                   :   std_logic_vector((RX_DATA_WIDTH-1) downto 0);
    signal  rx_data_r_track             :   std_logic_vector((RX_DATA_WIDTH-1) downto 0);
    signal  start_of_packet_detected_r  :   std_logic;    
    signal  track_data_r                :   std_logic;
    signal  track_data_r2               :   std_logic;
    signal  track_data_r3               :   std_logic;
    signal  rx_data_r2                  :   std_logic_vector((RX_DATA_WIDTH-1) downto 0);
    signal  rx_data_r3                  :   std_logic_vector((RX_DATA_WIDTH-1) downto 0);
    signal  rx_data_r4                  :   std_logic_vector((RX_DATA_WIDTH-1) downto 0);
    signal  rx_data_r5                  :   std_logic_vector((RX_DATA_WIDTH-1) downto 0);
    signal  rx_data_r6                  :   std_logic_vector((RX_DATA_WIDTH-1) downto 0);
    signal  rxctrl_r                    :   std_logic_vector((RXCTRL_WIDTH-1) downto 0);
    signal  rxctrl_r2                   :   std_logic_vector((RXCTRL_WIDTH-1) downto 0);
    signal  rxctrl_r3                   :   std_logic_vector((RXCTRL_WIDTH-1) downto 0);

    signal  rx_chanbond_seq_r           :   std_logic;
    signal  rx_chanbond_seq_r2          :   std_logic;
    signal  rx_chanbond_seq_r3          :   std_logic;
 
    signal  idle_slip_r                 :   std_logic;
    signal  slip_assert_r               :   std_logic;
    signal  wait_state_r                :   std_logic;
    signal  bit_align_r                 :   std_logic;
    signal  wait_before_slip_r          :   std_logic_vector(6 downto 0);
    signal  wait_before_init_r          :   std_logic_vector(6 downto 0);
 
    signal  sel                         :   std_logic_vector(1 downto 0);
 
    signal  rx_chanbond_reg_bitwise_or_i:   std_logic; 
 

--*********************************Wire Declarations***************************
   
    signal  bram_data_r                 :   std_logic_vector((RX_DATA_WIDTH-1) downto 0);
    signal  rx_data_ram_r               :   std_logic_vector(79 downto 0);
    signal  error_detected_c            :   std_logic;
    signal  input_to_chanbond_data_i    :   std_logic;
    signal  input_to_chanbond_reg_i     :   std_logic;
    signal  chanbondseq_in_data         :   std_logic;
    signal  rx_chanbond_reg             :   std_logic_vector((CHANBOND_SEQ_LEN-1) downto 0);
    signal  rxdata_or                   :   std_logic;
    signal  rxdata_r_or                 :   std_logic;
    signal  rxdata_r2_or                :   std_logic;
    signal  rxdata_r3_or                :   std_logic;
    signal  count_slip_complete_c       :   std_logic;
    signal  next_idle_slip_c            :   std_logic;
    signal  next_slip_assert_c          :   std_logic;
    signal  wait_state_c                :   std_logic;
    signal  rx_data_aligned             :   std_logic_vector((RX_DATA_WIDTH-1) downto 0);
    signal  next_begin_c                :   std_logic;
    signal  next_data_error_detected_c  :   std_logic;
    signal  next_track_data_c           :   std_logic;
    signal  start_of_packet_detected_c  :   std_logic;
    signal  rx_data_has_start_char_c    :   std_logic;
    signal  rx_data_matches_bram_c      :   std_logic;
    signal  tied_to_ground_i            :   std_logic;
    signal  tied_to_ground_vec_i        :   std_logic_vector(31 downto 0);
    signal  tied_to_vcc_i               :   std_logic;


--*********************************User Defined Attribute*****************************

    type RomType is array(0 to 511) of std_logic_vector(79 downto 0);
    type check_type is(
    ST_LINK_DOWN, ST_LINK_UP);
    
  signal sm_link : std_logic := '0';
  signal link_ctr : std_logic_vector(6 downto 0) := "0000000";

    impure function InitRomFromFile (RomFileName : in string) return RomType is

         FILE RomFile : text open read_mode is RomFileName;
         variable RomFileLine : line;
         variable ROM : RomType;
    begin
         for i in RomType'range loop
           readline (RomFile, RomFileLine);
           hread (RomFileLine, ROM(i));
         end loop;
         return ROM;
    end function;

    signal ROM : RomType := InitRomFromFile("gt_rom_init_rx.dat");


   function or_reduce(arg: std_logic_vector) return std_logic is
	variable result: std_logic;
    begin
	result := '0';
	for i in arg'range loop
	    result := result or arg(i);
	end loop;
        return result;
    end;

--*********************************Main Body of Code***************************
begin

    --_______________________  Static signal Assigments _______________________   

    tied_to_ground_i        <= '0';
    tied_to_ground_vec_i    <= (others=>'0');
    tied_to_vcc_i           <= '1';

    --___________ synchronizing the async reset for ease of timing simulation ________
    process( USER_CLK )
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            system_reset_r <= SYSTEM_RESET after DLY; 
            system_reset_r2 <= system_reset_r after DLY; 
        end if;
    end process; 

    process( USER_CLK )
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            reset_on_error_in_r <= RESET_ON_ERROR_IN after DLY; 
            reset_on_error_in_r2 <= reset_on_error_in_r after DLY; 
        end if;
    end process;    

    --______________________ Register RXDATA once to ease timing ______________   

    process( USER_CLK )
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            rx_data_r  <= RX_DATA_IN   after DLY;
            rx_data_r2 <= rx_data_r    after DLY;
        end if;
    end process;

    process( USER_CLK )
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            rxctrl_r   <= RXCTRL_IN   after DLY;
        end if;
    end process;
    --________________________________ State machine __________________________    
    
    
    -- State registers
    process( USER_CLK )
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            if(system_reset_r2 = '1') then
                begin_r                <=  '1' after DLY;
                track_data_r           <=  '0' after DLY;
                data_error_detected_r  <=  '0' after DLY;
            else
                begin_r                <=  next_begin_c after DLY;
                track_data_r           <=  next_track_data_c after DLY;
                data_error_detected_r  <=  next_data_error_detected_c after DLY;
            end if;
        end if;
    end process;

    -- Next state logic
    next_begin_c               <=   (begin_r and not start_of_packet_detected_r) or data_error_detected_r ;

    next_track_data_c          <=   (begin_r and start_of_packet_detected_r) or (track_data_r and not error_detected_r);
                                      
    next_data_error_detected_c <=   (track_data_r and error_detected_r);                               
        
    start_of_packet_detected_c <=   rx_data_has_start_char_c;

    process( USER_CLK )
    begin
    if(USER_CLK'event and USER_CLK = '1') then
        start_of_packet_detected_r    <=   start_of_packet_detected_c after DLY;
    end if;    
    end process;
    
    -- Registering for timing
    process( USER_CLK )
    begin
    if(USER_CLK'event and USER_CLK = '1') then
        track_data_r2    <=   track_data_r after DLY;
    end if;    
    end process;

    process( USER_CLK )
    begin
    if(USER_CLK'event and USER_CLK = '1') then
        track_data_r3    <=   track_data_r2 after DLY;
    end if;    
    end process;

    --______________________________ Capture incoming data ____________________    

    process( USER_CLK )
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            if(system_reset_r2 = '1') then 
                rx_data_r3      <=  (others => '0') after DLY;
            else
                if(sel = "01")  then
                    rx_data_r3  <=  rx_data_r((RX_DATA_WIDTH/2 - 1) downto 0) & rx_data_r2((RX_DATA_WIDTH-1) downto RX_DATA_WIDTH/2) after DLY;  
                else              
                    rx_data_r3  <=  rx_data_r2 after DLY;
                end if;    
            end if; 
        end if;
    end process;

    process( USER_CLK )
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            if(system_reset_r2 = '1') then 
                rx_data_r4      <=  (others => '0') after DLY;
                rx_data_r5      <=  (others => '0') after DLY;
                rx_data_r6      <=  (others => '0') after DLY;
                rx_data_r_track <=  (others => '0') after DLY;
            else
                rx_data_r4      <=  rx_data_r3 after DLY;
                rx_data_r5      <=  rx_data_r4 after DLY;
                rx_data_r6      <=  rx_data_r5 after DLY;
                rx_data_r_track <=  rx_data_r6 after DLY;
            end if;
        end if;    
    end process;

    process( USER_CLK )
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            if(system_reset_r2 = '1') then 
                rxctrl_r2      <=  (others => '0') after DLY;
                rxctrl_r3      <=  (others => '0') after DLY;
            else
                rxctrl_r2      <=  rxctrl_r  after DLY;
                rxctrl_r3      <=  rxctrl_r2 after DLY;
            end if;
        end if;    
    end process;

    rx_data_aligned <= rx_data_r3;

    -- ___________________________ Code for Channel bonding ____________________    
    -- code to prevent checking of clock correction sequences for the start of packet char
    process( USER_CLK )
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            rx_chanbond_seq_r    <=  RX_CHANBOND_SEQ_IN after DLY;
            rx_chanbond_seq_r2   <=  rx_chanbond_seq_r after DLY;
            rx_chanbond_seq_r3   <=  rx_chanbond_seq_r2 after DLY;
        end if;    
    end process;

    input_to_chanbond_reg_i  <= rx_chanbond_seq_r2;
    input_to_chanbond_data_i <= tied_to_ground_i;

   --______________ Code for Bit Slipping Logic______________
   
    process(rx_data_r)
    variable or_rxdata_r_var : std_logic;
    variable i             : std_logic;
    begin
        or_rxdata_r_var := '0';
        bit_wise_rxdata_r_or : for  i in 0 to (RX_DATA_WIDTH-1) loop
            or_rxdata_r_var :=  or_rxdata_r_var or rx_data_r(i);
        end loop;
        rxdata_r_or <= or_rxdata_r_var;
    end process;

    process(rx_data_r2)
    variable or_rxdata_r2_var : std_logic;
    variable i             : std_logic;
    begin
        or_rxdata_r2_var := '0';
        bit_wise_rxdata_r2_or : for  i in 0 to (RX_DATA_WIDTH-1) loop
            or_rxdata_r2_var :=  or_rxdata_r2_var or rx_data_r2(i);
        end loop;
        rxdata_r2_or <= or_rxdata_r2_var;
    end process;

    process(rx_data_r3)
    variable or_rxdata_r3_var : std_logic;
    variable i             : std_logic;
    begin
        or_rxdata_r3_var := '0';
        bit_wise_rxdata_r3_or : for  i in 0 to (RX_DATA_WIDTH-1) loop
            or_rxdata_r3_var :=  or_rxdata_r3_var or rx_data_r3(i);
        end loop;
        rxdata_r3_or <= or_rxdata_r3_var;
    end process;

    rxdata_or <= rxdata_r_or or rxdata_r2_or or rxdata_r3_or;

    -- State registers
    process( USER_CLK )
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            if( (system_reset_r2 = '1') or (wait_before_init_r(6) = '0') or (rxdata_or = '0') )then
                idle_slip_r            <=  '1' after DLY;
                slip_assert_r          <=  '0' after DLY;
                wait_state_r           <=  '0' after DLY;
            else
                idle_slip_r            <=  next_idle_slip_c   after DLY;
                slip_assert_r          <=  next_slip_assert_c after DLY;
                wait_state_r           <=  wait_state_c       after DLY;
            end if;
        end if;
    end process;
 
    -- Next state logic
    next_idle_slip_c           <=   (idle_slip_r and bit_align_r) or (wait_state_r and count_slip_complete_c) ;     

    next_slip_assert_c         <=   (idle_slip_r and (not bit_align_r));

    wait_state_c               <=   (slip_assert_r) or (wait_state_r and (not count_slip_complete_c)); 


    --_______ Counter for waiting clock cycles after RXSLIDE________
    process( USER_CLK )
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            if(wait_state_r = '0') then
               wait_before_slip_r  <=  "0000000" after DLY;
            else
               wait_before_slip_r  <=  wait_before_slip_r + '1' after DLY;
            end if;
        end if;
    end process;

    --_______ Counter for waiting clock cycles before starting RXSLIDE operation________
    --_______ Wait for 64 clock cycles to see if the RXDATA is already byte aligned. If not, start RXSLIDE operation
    process( USER_CLK )
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            if( (system_reset_r2 = '1') or (rxdata_or = '0') ) then
               wait_before_init_r  <=  "0000000" after DLY;
            elsif(wait_before_init_r(6) = '0') then 
               wait_before_init_r  <=  wait_before_init_r + '1' after DLY;
            end if;
        end if;
    end process;

    count_slip_complete_c <= wait_before_slip_r(6);

    process( USER_CLK )
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            if( (system_reset_r2 = '1') or (rxdata_or = '0') ) then
                  bit_align_r  <=  '0'  after DLY;
            else 
                if( ((rx_data_r(7 downto 0) & rx_data_r2(15 downto 8)) = START_OF_PACKET_CHAR) or (rx_data_r(15 downto 0) = START_OF_PACKET_CHAR) ) then
 
                     bit_align_r   <=   '1'  after DLY;
                
                end if;
            end if;
        end if;
    end process;


    -- In 2 Byte scenario, when align_comma_word=1, Comma can appear on any of the two bytes
    -- The comma is moved to the lower byte so that error checking can start
    process( USER_CLK )
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            if((reset_on_error_in_r2='1') or (system_reset_r2='1')) then 
                sel <= "00";
            elsif ((begin_r= '1') and (rx_chanbond_seq_r = '0')) then
             -- if Comma appears on BYTE0 ..
                if((rx_data_r((RX_DATA_WIDTH/2 - 1) downto 0) = START_OF_PACKET_CHAR(7 downto 0))  and (rxctrl_r(0) = '1'))then
                    sel <= "00";
             -- if Comma appears on BYTE1 ..     
                elsif((rx_data_r((RX_DATA_WIDTH-1) downto RX_DATA_WIDTH/2) = START_OF_PACKET_CHAR(7 downto 0))  and (rxctrl_r(1) = '1'))then
                    sel <= "01";
                end if;
            end if;
        end if;
    end process;
    --___________________________ Code for Channel bonding ____________________    
    -- code to prevent checking of clock correction sequences for the start of packet char
    register_chan_seq: for i in 0 to (CHANBOND_SEQ_LEN-1) generate
        case_i_equal_to_0: if (i=0) generate 
            rx_chanbond_reg_0 : FD port map (Q => rx_chanbond_reg(i),D => input_to_chanbond_reg_i,C => USER_CLK);
        end generate case_i_equal_to_0;
        case_i_greater_than_0: if (i>0) generate 
            rx_chanbond_reg_i :FD port map (Q => rx_chanbond_reg(i),D => rx_chanbond_reg(i-1),C => USER_CLK);
        end generate case_i_greater_than_0;
    end generate register_chan_seq;
    
    chanbondseq_in_data <= input_to_chanbond_data_i or rx_chanbond_reg_bitwise_or_i;

    process(rx_chanbond_reg)
    variable rx_chanbond_var : std_logic;
    variable i               : std_logic;
    begin
        rx_chanbond_var := '0';
        bit_wise_or : for  i in 0 to (CHANBOND_SEQ_LEN-1) loop
            rx_chanbond_var :=  rx_chanbond_var or rx_chanbond_reg(i);
        end loop;
        rx_chanbond_reg_bitwise_or_i <= rx_chanbond_var;
    end process;

    rx_data_has_start_char_c <= '1' when ((rx_data_aligned(7 downto 0) = START_OF_PACKET_CHAR(7 downto 0)) and (chanbondseq_in_data='0') and (or_reduce(rxctrl_r3)='1')) else '0';


    --_____________________________ Assign output ports _______________________    


    --TRACK_DATA_OUT      <=  track_data_r;  

    RX_SLIDE            <=  slip_assert_r;

    -- Drive the enpcommaalign port of the gt for alignment
    process( USER_CLK )
    begin
    if(USER_CLK'event and USER_CLK = '1') then
        if(system_reset_r2 = '1') then 
            RXENPCOMMADET_OUT   <= '0' after DLY;
        else              
            RXENPCOMMADET_OUT   <= '1' after DLY;
        end if;
    end if;    
    end process;

    -- Drive the enmcommaalign port of the gt for alignment
    process( USER_CLK )
    begin
    if(USER_CLK'event and USER_CLK = '1') then
        if(system_reset_r2 = '1') then 
            RXENMCOMMADET_OUT   <= '0' after DLY;
        else              
            RXENMCOMMADET_OUT   <= '1' after DLY;
        end if;
    end if;    
    end process;

    INC_OUT            <=  start_of_packet_detected_c;   

    PATTERN_MATCHB_OUT <=  data_error_detected_r;

    -- Drive the enchansync port of the mgt for channel bonding
    process( USER_CLK )
    begin
    if(USER_CLK'event and USER_CLK = '1') then
        if(system_reset_r2 = '1') then 
            RX_ENCHAN_SYNC_OUT   <= '0' after DLY;
        else              
            RX_ENCHAN_SYNC_OUT   <= '1' after DLY;
        end if;
    end if;    
    end process;

    --___________________________ Check incoming data for errors ______________
         
    
    --An error is detected when data read for the BRAM does not match the incoming data

    rx_data_matches_bram_c <= '0' when (rx_data_r_track /= bram_data_r) else '1';

    error_detected_c    <=   track_data_r3 and not rx_data_matches_bram_c;   
    
    --We register the error_detected signal for use with the error counter logic
    process( USER_CLK )
    begin
    if(USER_CLK'event and USER_CLK = '1') then
        if(not(track_data_r = '1')) then 
            error_detected_r    <= '0' after DLY;
        else
            error_detected_r    <=  error_detected_c after DLY;
        end if;
    end if;    
    end process;

    --We count the total number of errors we detect. By keeping a count we make it less likely that we will miss
    --errors we did not directly observe. This counter must be reset when it reaches its max value
    process ( USER_CLK )
    begin
    if( USER_CLK'event and USER_CLK = '1') then
        if(system_reset_r2='1') then
            error_count_r       <=  (others => '0') after DLY;
        elsif(error_detected_r = '1') then
            error_count_r       <=  error_count_r + 1 after DLY;
        end if;
    end if;
    end process;
            
    --Here we connect the lower 8 bits of the count (the MSbit is used only to check when the counter reaches
    --max value) to the module output
    ERROR_COUNT_OUT     <=   std_logic_vector(error_count_r(7 downto 0));



process(USER_CLK)
  begin
    if( USER_CLK'event and USER_CLK = '1') then
       if(track_data_r='0') then
             sm_link  <= '0';
       else
    case sm_link is
      -- The link is considered to be down when the link counter initially has a value less than 67. When the link is
      -- down, the counter is incremented on each cycle where all PRBS bits match, but reset whenever any PRBS mismatch
      -- occurs. When the link counter reaches 67, transition to the link up state.
       when '0' =>
        if (error_detected_r = '1') then
          link_ctr <= (others => '0');
        else 
          if (link_ctr < "1000011") then
            link_ctr <= link_ctr + '1';
          else
            sm_link <= '1';
        end if;
      end if;

      -- When the link is up, the link counter is decreased by 34 whenever any PRBS mismatch occurs, but is increased by
      -- only 1 on each cycle where all PRBS bits match, up to its saturation point of 67. If the link counter reaches
      -- 0 (including rollover protection), transition to the link down state.
       when '1' => 
        if (error_detected_r = '1') then
          if (link_ctr > "0100001") then
            link_ctr <= link_ctr - "0100010";
            if (link_ctr = "0100010") then
              sm_link  <= '0';
            end if;
          else 
            link_ctr <= (others => '0');
            sm_link  <= '0';
          end if;
        else 
          if (link_ctr < "1000011") then
            link_ctr <= link_ctr + '1';
        end if;
      end if;
       when OTHERS =>
            sm_link  <= '0';
    end case;
  end if;
  end if;
 end process; 

   TRACK_DATA_OUT <= sm_link;

    --____________________________ Counter to read from BRAM __________________________    
    process( USER_CLK )
    begin
    if(USER_CLK'event and USER_CLK = '1') then
        if((system_reset_r2='1') or (read_counter_i = (WORDS_IN_BRAM-1)))  then
            read_counter_i   <=  (others => '0') after DLY;
        elsif(((start_of_packet_detected_r and not track_data_r)='1')) then
            read_counter_i   <=  "0000000000" after DLY;
        else read_counter_i  <=  read_counter_i + 1 after DLY;
        end if;
    end if;
    end process;

    --________________________________ BRAM Inference Logic _____________________________    

--Array slice from dat file to compare against receive data
datapath_80 : if(RX_DATA_WIDTH = 80) generate
begin
    bram_data_r         <= rx_data_ram_r((RX_DATA_WIDTH-1) downto 0);
end generate datapath_80;

datapath_16_20_32_40_64 : if((RX_DATA_WIDTH = 16) or (RX_DATA_WIDTH = 20) or (RX_DATA_WIDTH = 32) or (RX_DATA_WIDTH = 40) or (RX_DATA_WIDTH = 64)) generate
begin
    bram_data_r         <= rx_data_ram_r((16+RX_DATA_WIDTH-1) downto 16);
end generate datapath_16_20_32_40_64;

    read_counter_conv   <= std_logic_vector(read_counter_i);

    process (USER_CLK)
    begin
       if(USER_CLK'event and USER_CLK='1') then
         rx_data_ram_r <= ROM(conv_integer(read_counter_conv)) after DLY;
       end if;
    end process;
    
    
end RTL;           

